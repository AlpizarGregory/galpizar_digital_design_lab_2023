module mux_dibujar(

	input logic line,
	input logic [23:0]rgb0,rgb1,rgb2,rgb3,rgb4,rgb5,rgb6,rgb7,rgb8,rgb9,rgb10,rgb11,rgb12,rgb13,rgb14,rgb15,rgb16,rgb17,rgb18,rgb19,rgb20,rgb21,rgb22,rgb23,rgb24,rgb25,rgb26,rgb27,rgb28,rgb29,rgb30,rgb31,rgb32,rgb33,rgb34,rgb35,rgb36,rgb37,rgb38,rgb39,rgb40,rgb41,rgb42,rgb43,rgb44,rgb45,rgb46,rgb47,rgb48,rgb49,rgb50,rgb51,rgb52,rgb53,rgb54,rgb55,rgb56,rgb57,rgb58,rgb59,rgb60,rgb61,rgb62,rgb63,
	input logic pos0,pos1,pos2,pos3,pos4,pos5,pos6,pos7,pos8,pos9,pos10,pos11,pos12,pos13,pos14,pos15,pos16,pos17,pos18,pos19,pos20,pos21,pos22,pos23,pos24,pos25,pos26,pos27,pos28,pos29,pos30,pos31,pos32,pos33,pos34,pos35,pos36,pos37,pos38,pos39,pos40,pos41,pos42,pos43,pos44,pos45,pos46,pos47,pos48,pos49,pos50,pos51,pos52,pos53,pos54,pos55,pos56,pos57,pos58,pos59,pos60,pos61,pos62,pos63,
	input logic win,lose,
	output logic [7:0]r,g,b

);

	logic[23:0]out_rgb;
	
	always_comb begin   

		case({line,pos0,pos1,pos2,pos3,pos4,pos5,pos6,pos7,pos8,pos9,pos10,pos11,pos12,pos13,pos14,pos15,pos16,pos17,pos18,pos19,pos20,pos21,pos22,pos23,pos24,pos25,pos26,pos27,pos28,pos29,pos30,pos31,pos32,pos33,pos34,pos35,pos36,pos37,pos38,pos39,pos40,pos41,pos42,pos43,pos44,pos45,pos46,pos47,pos48,pos49,pos50,pos51,pos52,pos53,pos54,pos55,pos56,pos57,pos58,pos59,pos60,pos61,pos62,pos63,win,lose})
		
			67'b0000000000000000000000000000000000000000000000000000000000000000010 : out_rgb <= 24'h00FF00;
			67'b0000000000000000000000000000000000000000000000000000000000000000001 : out_rgb <= 24'hFF0000;
			67'b0000000000000000000000000000000000000000000000000000000000000000000 : out_rgb <= 24'h000000;
			67'b1000000000000000000000000000000000000000000000000000000000000000000 : out_rgb <= 24'hffffff;
			67'b0100000000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb0;
			67'b0010000000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb1;
			67'b0001000000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb2;
			67'b0000100000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb3;
			67'b0000010000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb4;
			67'b0000001000000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb5;
			67'b0000000100000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb6;
			67'b0000000010000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb7;
			67'b0000000001000000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb8;
			67'b0000000000100000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb9;
			67'b0000000000010000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb10;
			67'b0000000000001000000000000000000000000000000000000000000000000000000 : out_rgb <= rgb11;
			67'b0000000000000100000000000000000000000000000000000000000000000000000 : out_rgb <= rgb12;
			67'b0000000000000010000000000000000000000000000000000000000000000000000 : out_rgb <= rgb13;
			67'b0000000000000001000000000000000000000000000000000000000000000000000 : out_rgb <= rgb14;
			67'b0000000000000000100000000000000000000000000000000000000000000000000 : out_rgb <= rgb15;
			67'b0000000000000000010000000000000000000000000000000000000000000000000 : out_rgb <= rgb16;
			67'b0000000000000000001000000000000000000000000000000000000000000000000 : out_rgb <= rgb17;
			67'b0000000000000000000100000000000000000000000000000000000000000000000 : out_rgb <= rgb18;
			67'b0000000000000000000010000000000000000000000000000000000000000000000 : out_rgb <= rgb19;
			67'b0000000000000000000001000000000000000000000000000000000000000000000 : out_rgb <= rgb20;
			67'b0000000000000000000000100000000000000000000000000000000000000000000 : out_rgb <= rgb21;
			67'b0000000000000000000000010000000000000000000000000000000000000000000 : out_rgb <= rgb22;
			67'b0000000000000000000000001000000000000000000000000000000000000000000 : out_rgb <= rgb23;
			67'b0000000000000000000000000100000000000000000000000000000000000000000 : out_rgb <= rgb24;
			67'b0000000000000000000000000010000000000000000000000000000000000000000 : out_rgb <= rgb25;
			67'b0000000000000000000000000001000000000000000000000000000000000000000 : out_rgb <= rgb26;
			67'b0000000000000000000000000000100000000000000000000000000000000000000 : out_rgb <= rgb27;
			67'b0000000000000000000000000000010000000000000000000000000000000000000 : out_rgb <= rgb28;
			67'b0000000000000000000000000000001000000000000000000000000000000000000 : out_rgb <= rgb29;
			67'b0000000000000000000000000000000100000000000000000000000000000000000 : out_rgb <= rgb30;
			67'b0000000000000000000000000000000010000000000000000000000000000000000 : out_rgb <= rgb31;
			67'b0000000000000000000000000000000001000000000000000000000000000000000 : out_rgb <= rgb32;
			67'b0000000000000000000000000000000000100000000000000000000000000000000 : out_rgb <= rgb33;
			67'b0000000000000000000000000000000000010000000000000000000000000000000 : out_rgb <= rgb34;
			67'b0000000000000000000000000000000000001000000000000000000000000000000 : out_rgb <= rgb35;
			67'b0000000000000000000000000000000000000100000000000000000000000000000 : out_rgb <= rgb36;
			67'b0000000000000000000000000000000000000010000000000000000000000000000 : out_rgb <= rgb37;
			67'b0000000000000000000000000000000000000001000000000000000000000000000 : out_rgb <= rgb38;
			67'b0000000000000000000000000000000000000000100000000000000000000000000 : out_rgb <= rgb39;
			67'b0000000000000000000000000000000000000000010000000000000000000000000 : out_rgb <= rgb40;
			67'b0000000000000000000000000000000000000000001000000000000000000000000 : out_rgb <= rgb41;
			67'b0000000000000000000000000000000000000000000100000000000000000000000 : out_rgb <= rgb42;
			67'b0000000000000000000000000000000000000000000010000000000000000000000 : out_rgb <= rgb43;
			67'b0000000000000000000000000000000000000000000001000000000000000000000 : out_rgb <= rgb44;
			67'b0000000000000000000000000000000000000000000000100000000000000000000 : out_rgb <= rgb45;
			67'b0000000000000000000000000000000000000000000000010000000000000000000 : out_rgb <= rgb46;
			67'b0000000000000000000000000000000000000000000000001000000000000000000 : out_rgb <= rgb47;
			67'b0000000000000000000000000000000000000000000000000100000000000000000 : out_rgb <= rgb48;
			67'b0000000000000000000000000000000000000000000000000010000000000000000 : out_rgb <= rgb49;
			67'b0000000000000000000000000000000000000000000000000001000000000000000 : out_rgb <= rgb50;
			67'b0000000000000000000000000000000000000000000000000000100000000000000 : out_rgb <= rgb51;
			67'b0000000000000000000000000000000000000000000000000000010000000000000 : out_rgb <= rgb52;
			67'b0000000000000000000000000000000000000000000000000000001000000000000 : out_rgb <= rgb53;
			67'b0000000000000000000000000000000000000000000000000000000100000000000 : out_rgb <= rgb54;
			67'b0000000000000000000000000000000000000000000000000000000010000000000 : out_rgb <= rgb55;
			67'b0000000000000000000000000000000000000000000000000000000001000000000 : out_rgb <= rgb56;
			67'b0000000000000000000000000000000000000000000000000000000000100000000 : out_rgb <= rgb57;
			67'b0000000000000000000000000000000000000000000000000000000000010000000 : out_rgb <= rgb58;
			67'b0000000000000000000000000000000000000000000000000000000000001000000 : out_rgb <= rgb59;
			67'b0000000000000000000000000000000000000000000000000000000000000100000 : out_rgb <= rgb60;
			67'b0000000000000000000000000000000000000000000000000000000000000010000 : out_rgb <= rgb61;
			67'b0000000000000000000000000000000000000000000000000000000000000001000 : out_rgb <= rgb62;
			67'b0000000000000000000000000000000000000000000000000000000000000000100 : out_rgb <= rgb63;
		

				 // 0    1    2    3     4   5    6    7    8    9    A     B     C     D     E     F     G
			//case ({line,pos0,pos1,pos2,pos3,pos4,pos5,pos6,pos7,pos8,pos9,pos10,pos11,pos12,pos13,pos14,pos15,win,lose})
			//
			//19'b0000000000000000000 : out_rgb     <= 24'h000000;
			//19'b1000000000000000000 : out_rgb     <= 24'hffffff;
			//19'b0100000000000000000 : out_rgb     <= rgb0;
			//19'b0010000000000000000 : out_rgb     <= rgb1;
			//19'b0001000000000000000 : out_rgb     <= rgb2;
			//19'b0000100000000000000 : out_rgb     <= rgb3;
			//19'b0000010000000000000 : out_rgb     <= rgb4;
			//19'b0000001000000000000 : out_rgb     <= rgb5;
			//19'b0000000100000000000 : out_rgb     <= rgb6;
			//19'b0000000010000000000 : out_rgb     <= rgb7;
			//19'b0000000001000000000 : out_rgb     <= rgb8;
			//19'b0000000000100000000 : out_rgb     <= rgb9;
			//19'b0000000000010000000 : out_rgb     <= rgb10;
			//19'b0000000000001000000 : out_rgb     <= rgb11;
			//19'b0000000000000100000 : out_rgb     <= rgb12;
			//19'b0000000000000010000 : out_rgb     <= rgb13;
			//19'b0000000000000001000 : out_rgb     <= rgb14;
			//19'b0000000000000000100 : out_rgb     <= rgb15;
			//  //0123456789ABCDEFG
			//
			////Casos win/lose
			//19'b1000000000000000010 : out_rgb     <= 24'b000000000000000011111111;
			//19'b1000000000000000001 : out_rgb     <= 24'b111111110000000000000000;
			
			default  : out_rgb <= 24'hA7A200;
			
		endcase
	end
		
	assign r = out_rgb[23:16];
	assign g = out_rgb[15:8];
	assign b = out_rgb[7:0];
	
endmodule
module CheckPos(input logic [9:0] hs,vs,
				output logic [63:0]pos);
		//logic paint;		  
		//for (i = 0; i < 64; i++) begin
		//	paint = 
		//end

		//assign pos[0]  = ((5   < hs)&(151 > hs)&(5   < vs)&(110 > vs))? 1:0;
		//assign pos[1]  = ((171 < hs)&(311 > hs)&(5   < vs)&(110 > vs))? 1:0;
		//assign pos[2]  = ((331 < hs)&(471 > hs)&(5   < vs)&(110 > vs))? 1:0;
		//assign pos[3]  = ((491 < hs)&(631 > hs)&(5   < vs)&(110 > vs))? 1:0;
		//assign pos[4]  = ((5   < hs)&(151 > hs)&(130 < vs)&(230 > vs))? 1:0;
		//assign pos[5]  = ((171 < hs)&(311 > hs)&(130 < vs)&(230 > vs))? 1:0;
		//assign pos[6]  = ((331 < hs)&(471 > hs)&(130 < vs)&(230 > vs))? 1:0;
		//assign pos[7]  = ((491 < hs)&(631 > hs)&(130 < vs)&(230 > vs))? 1:0;
		//assign pos[8]  = ((5   < hs)&(151 > hs)&(250 < vs)&(350 > vs))? 1:0;
		//assign pos[9]  = ((171 < hs)&(311 > hs)&(250 < vs)&(350 > vs))? 1:0;
		//assign pos[10] = ((331 < hs)&(471 > hs)&(250 < vs)&(350 > vs))? 1:0;
		//assign pos[11] = ((491 < hs)&(631 > hs)&(250 < vs)&(350 > vs))? 1:0;
		//assign pos[12] = ((5   < hs)&(151 > hs)&(375 < vs)&(475 > vs))? 1:0;
		//assign pos[13] = ((171 < hs)&(311 > hs)&(375 < vs)&(475 > vs))? 1:0;
		//assign pos[14] = ((331 < hs)&(471 > hs)&(375 < vs)&(475 > vs))? 1:0;
		//assign pos[15] = ((491 < hs)&(631 > hs)&(375 < vs)&(475 > vs))? 1:0;
		
endmodule
module countdownNbits7seg
	#(parameter Nbits = 4)
		(input logic clk, reset, input logic [Nbits-1:0] first,
		output logic [13:0] seg);
	
	logic [Nbits-1:0] current;
	
	// asynchronous reset
	always @ (posedge clk, posedge reset)
		if (reset) current <= first;
		else current <= current - 1;
		//else current <= current;
	
	//always @ (negedge subtrac)
	//	if (subtrac) current <= current - 1;
	
	always @ (posedge clk)
		case(current)
			//			Two 7 segment display (HEX)
			
			'b000000: seg = 14'b1111111_0000001;
			'b000001: seg = 14'b1111111_1001111;
			'b000010: seg = 14'b1111111_0010010;
			'b000011: seg = 14'b1111111_0000110;
			'b000100: seg = 14'b1111111_1001100;
			'b000101: seg = 14'b1111111_0100100;
			'b000110: seg = 14'b1111111_0100000;
			'b000111: seg = 14'b1111111_0001111;
			'b001000: seg = 14'b1111111_0000000;
			'b001001: seg = 14'b1111111_0000100;
			//	
			'b001010: seg = 14'b1001111_0000001;
			'b001011: seg = 14'b1001111_1001111;
			'b001100: seg = 14'b1001111_0010010;
			'b001101: seg = 14'b1001111_0000110;
			'b001110: seg = 14'b1001111_1001100;
			'b001111: seg = 14'b1001111_0100100;
			'b010000: seg = 14'b1001111_0100000;
			'b010001: seg = 14'b1001111_0001111;
			'b010010: seg = 14'b1001111_0000000;
			'b010011: seg = 14'b1001111_0000100;
			//
			'b010100: seg = 14'b0010010_0000001;
			'b010101: seg = 14'b0010010_1001111;
			'b010110: seg = 14'b0010010_0010010;
			'b010111: seg = 14'b0010010_0000110;
			'b011000: seg = 14'b0010010_1001100;
			'b011001: seg = 14'b0010010_0100100;
			'b011010: seg = 14'b0010010_0100000;
			'b011011: seg = 14'b0010010_0001111;
			'b011100: seg = 14'b0010010_0000000;
			'b011101: seg = 14'b0010010_0000100;
			//
			'b011110: seg = 14'b0000110_0000001;
			'b011111: seg = 14'b0000110_1001111;
			'b100000: seg = 14'b0000110_0010010;
			'b100001: seg = 14'b0000110_0000110;
			'b100010: seg = 14'b0000110_1001100;
			'b100011: seg = 14'b0000110_0100100;
			'b100100: seg = 14'b0000110_0100000;
			'b100101: seg = 14'b0000110_0001111;
			'b100110: seg = 14'b0000110_0000000;
			'b100111: seg = 14'b0000110_0000100;
			//
			'b101000: seg = 14'b1001100_0000001;
			'b101001: seg = 14'b1001100_1001111;
			'b101010: seg = 14'b1001100_0010010;
			'b101011: seg = 14'b1001100_0000110;
			'b101100: seg = 14'b1001100_1001100;
			'b101101: seg = 14'b1001100_0100100;
			'b101110: seg = 14'b1001100_0100000;
			'b101111: seg = 14'b1001100_0001111;
			'b110000: seg = 14'b1001100_0000000;
			'b110001: seg = 14'b1001100_0000100;
			//
			'b110010: seg = 14'b0100100_0000001;
			'b110011: seg = 14'b0100100_1001111;
			'b110100: seg = 14'b0100100_0010010;
			'b110101: seg = 14'b0100100_0000110;
			'b110110: seg = 14'b0100100_1001100;
			'b110111: seg = 14'b0100100_0100100;
			'b111000: seg = 14'b0100100_0100000;
			'b111001: seg = 14'b0100100_0001111;
			'b111010: seg = 14'b0100100_0000000;
			'b111011: seg = 14'b0100100_0000100;
			//
			'b111100: seg = 14'b0100000_0000001;
			'b111101: seg = 14'b0100000_1001111;
			'b111110: seg = 14'b0100000_0010010;
			'b111111: seg = 14'b0100000_0000110;
			default: seg = 14'b1111111_1111111;
			
		endcase
		
		

	
endmodule